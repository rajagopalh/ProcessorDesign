
module booth_encoder(y, x1_b, x2_b, Z, Neg); 
   



endmodule // booth_encoder

module booth_decoder(x, Neg, x1_b, x2_b, Z, PP);

endmodule // booth_decoder